`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 05/27/2019 07:00:37 AM
// Design Name:
// Module Name: tb
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

typedef struct packed {
    logic ap_clk;
    logic ap_rst;
    logic ap_start;
    logic ap_done;
    logic ap_idle;
    logic ap_ready;
} ap_ctrl;


typedef struct packed {
    logic tValid;
    logic [63:0] tData;
    logic [7:0] tUser;
    logic tLast;
} linkmastertype;

typedef struct packed {
    bit tReady;
} linkslavetype;

typedef struct {
    linkmastertype master;
    linkslavetype slave;
} axis;


function string wp_split(input int offset, string str, output int cnt);
    int i = 0;

    // Skip any existing whitespaces
    do begin
        if (str[offset] != " " && str[offset] != "\t") break;
    end while (++offset < str.len());

    if (offset == str.len()) begin
        cnt = 0;
        return "";
    end

    for (i = offset; i < str.len(); i++) begin
        if (str[i] == " " || str[i] == "\t") break;
    end

    cnt = i;
    return str.substr(offset,i-1);
endfunction

module tb ();
    // Parameters are set externally
    // With ruckus this is done by setting the SIM_PARAMETERS variable, for example:
    // make xsim SIM_PARAMETERS="tv_in=tv_in.txt tv_out=tv_out.txt"
    parameter tv_in="";
    parameter tv_out="";
    parameter tv_ref=""; // Not yet supported

    const string tv_in_str = tv_in;
    const string tv_out_str = tv_out;
    const string tv_ref_str = tv_ref;

    // Clock and reset signal declaration
    bit clk = 0;
    bit ready = 0;
    bit done = 0;

    ap_ctrl ctrl;           // HLS handshake signaling
    axis link_in[0:23];     // All AXI-stream inputs
    axis link_out[0:23];    // All AXI-stream outputs

    // Clock generation
    always #5 clk = ~clk;
    assign ctrl.ap_clk = clk;

    int fdr = 0, fdw = 0, fdref = 0;

    initial begin
        if (tv_in_str.len() == 0) $error("tv_in needs to be set");

        fdr = $fopen(tv_in_str, "r");
        if (fdr == 0) begin
            $error("Unable to open input file: %s", tv_in_str);
            $finish;
        end


        if (tv_out_str.len() == 0) begin
            $warning("tv_out isn't set, no output results will be written!");
        end else begin
            fdw = $fopen(tv_out_str, "w");
            if (fdw == 0) $error("Unable to open output file: %s", tv_out_str);

            $fwrite(fdw, "# Link output vector file from firmware RTL\n\n");
            // TODO: Work on the timestamp
            //$fdisplay(fdw, "# Generated by APx Gen2 testbench on %t", $timeformat(-9, 2, " ns", 20));
        end

        for (int i = 0; i < 24; i++) begin
            link_in[i].master.tValid = 0;
            link_in[i].master.tLast = 0;

            link_out[i].slave.tReady = 1;
        end

        // Reset and start logic
        ctrl.ap_rst = 1;
        ctrl.ap_start = 0;
        #25
        ctrl.ap_rst = 0;
        for (int i = 0; i < 3; i++) @(posedge clk);
        ready = 1;

        // Wait for done flag to be set
        @(posedge done);

        // Let the HLS block process the rest of the data
        // TODO: Put it as a parameter? clock count maybe?
        #1000

        $fclose(fdr);
        $fclose(fdw);
    end

    int cycle = 0;
    int linenr = 0;

    always @ (posedge clk) begin
        if (ready) cycle++;

        if (ready && !done) begin
            string line;
            int eof = 0;

            ctrl.ap_start = 1;

            while (1) begin
                linenr++;

                eof = $feof(fdr);
                if (eof) break;

                $fgets(line, fdr);

                // Skip empty lines and comments
                if ((line.len() >= 1) && (line[0] != "#") && ((line[0] >= " ") && (line[0] <= "~"))) break;
            end

            if (!eof) begin
                int offset = 0;

                string id = wp_split(offset, line, offset);
                //$display("id=%s", id);
                //$display("char=%d", line[0]);

                for (int i = 0; i < 24; i++) begin
                    string user = wp_split(offset, line, offset);
                    string data = wp_split(offset, line, offset);

                    if (user[0] == "-" && data[0] == "-") begin
                        // Skip AXI write
                        link_in[i].master.tUser = {8{1'bX}};
                        link_in[i].master.tData = {64{1'bX}};
                        link_in[i].master.tValid = 0;
                        link_in[i].master.tLast = 0;
                    end else begin
                        //$display("user(%d)=%s", i, user);
                        //$display("data(%d)=%s", i, data);

                        if (link_in[i].slave.tReady == 0) begin
                            $warning("tReady for link %0d in data cycle %0d isn't set!", i, cycle);
                        end

                        if (!$sscanf(user, "0x%2x", link_in[i].master.tUser) ||
                            !$sscanf(data, "0x%16x", link_in[i].master.tData)) begin
                            $error("Cannot parse link %0d at line %0d", i, linenr);
                        end

                        link_in[i].master.tValid = 1;
                        link_in[i].master.tLast = 1;
                    end

                end
            end else begin
                done = 1;
            end
        end

        if (done) begin
            // When the test vector is done we still send data so the HLS
            // block can process the rest of the data
            for (int i = 0; i < 24; i++) begin
                link_in[i].master.tUser = {8{1'bX}};
                link_in[i].master.tData = {64{1'bX}};
                link_in[i].master.tValid = 1;
                link_in[i].master.tLast = 1;
            end
        end
    end

    always @ (posedge clk) begin
        // Only write output if tv_out is defined
        if (ready && fdw) begin
            $fwrite(fdw, "%3d  ", cycle);

            for (int i = 0; i < 24; i++) begin
                if (link_out[i].master.tValid) begin
                    $fwrite(fdw, "0x%2x ", link_out[i].master.tUser);
                    $fwrite(fdw, "0x%16x  ", link_out[i].master.tData);
                end else begin
                    $fwrite(fdw, "-    ");
                    $fwrite(fdw, "-                   ");
                end
            end

            $fwrite(fdw, "\n");
        end
    end

    algo_top_sim_wrapper DUT (
        .ap_clk(ctrl.ap_clk),
        .ap_rst(ctrl.ap_rst),
        .ap_start(ctrl.ap_start),
        .ap_done(ctrl.ap_done),
        .ap_idle(ctrl.ap_idle),
        .ap_ready(ctrl.ap_ready),
        .link_in_master_0_tvalid(link_in[0].master.tValid),
        .link_in_master_0_tdata(link_in[0].master.tData),
        .link_in_master_0_tuser(link_in[0].master.tUser),
        .link_in_master_0_tlast(link_in[0].master.tLast),
        .link_in_slave_0_tready(link_in[0].slave.tReady),
        .link_in_master_1_tvalid(link_in[1].master.tValid),
        .link_in_master_1_tdata(link_in[1].master.tData),
        .link_in_master_1_tuser(link_in[1].master.tUser),
        .link_in_master_1_tlast(link_in[1].master.tLast),
        .link_in_slave_1_tready(link_in[1].slave.tReady),
        .link_in_master_2_tvalid(link_in[2].master.tValid),
        .link_in_master_2_tdata(link_in[2].master.tData),
        .link_in_master_2_tuser(link_in[2].master.tUser),
        .link_in_master_2_tlast(link_in[2].master.tLast),
        .link_in_slave_2_tready(link_in[2].slave.tReady),
        .link_in_master_3_tvalid(link_in[3].master.tValid),
        .link_in_master_3_tdata(link_in[3].master.tData),
        .link_in_master_3_tuser(link_in[3].master.tUser),
        .link_in_master_3_tlast(link_in[3].master.tLast),
        .link_in_slave_3_tready(link_in[3].slave.tReady),
        .link_in_master_4_tvalid(link_in[4].master.tValid),
        .link_in_master_4_tdata(link_in[4].master.tData),
        .link_in_master_4_tuser(link_in[4].master.tUser),
        .link_in_master_4_tlast(link_in[4].master.tLast),
        .link_in_slave_4_tready(link_in[4].slave.tReady),
        .link_in_master_5_tvalid(link_in[5].master.tValid),
        .link_in_master_5_tdata(link_in[5].master.tData),
        .link_in_master_5_tuser(link_in[5].master.tUser),
        .link_in_master_5_tlast(link_in[5].master.tLast),
        .link_in_slave_5_tready(link_in[5].slave.tReady),
        .link_in_master_6_tvalid(link_in[6].master.tValid),
        .link_in_master_6_tdata(link_in[6].master.tData),
        .link_in_master_6_tuser(link_in[6].master.tUser),
        .link_in_master_6_tlast(link_in[6].master.tLast),
        .link_in_slave_6_tready(link_in[6].slave.tReady),
        .link_in_master_7_tvalid(link_in[7].master.tValid),
        .link_in_master_7_tdata(link_in[7].master.tData),
        .link_in_master_7_tuser(link_in[7].master.tUser),
        .link_in_master_7_tlast(link_in[7].master.tLast),
        .link_in_slave_7_tready(link_in[7].slave.tReady),
        .link_in_master_8_tvalid(link_in[8].master.tValid),
        .link_in_master_8_tdata(link_in[8].master.tData),
        .link_in_master_8_tuser(link_in[8].master.tUser),
        .link_in_master_8_tlast(link_in[8].master.tLast),
        .link_in_slave_8_tready(link_in[8].slave.tReady),
        .link_in_master_9_tvalid(link_in[9].master.tValid),
        .link_in_master_9_tdata(link_in[9].master.tData),
        .link_in_master_9_tuser(link_in[9].master.tUser),
        .link_in_master_9_tlast(link_in[9].master.tLast),
        .link_in_slave_9_tready(link_in[9].slave.tReady),
        .link_in_master_10_tvalid(link_in[10].master.tValid),
        .link_in_master_10_tdata(link_in[10].master.tData),
        .link_in_master_10_tuser(link_in[10].master.tUser),
        .link_in_master_10_tlast(link_in[10].master.tLast),
        .link_in_slave_10_tready(link_in[10].slave.tReady),
        .link_in_master_11_tvalid(link_in[11].master.tValid),
        .link_in_master_11_tdata(link_in[11].master.tData),
        .link_in_master_11_tuser(link_in[11].master.tUser),
        .link_in_master_11_tlast(link_in[11].master.tLast),
        .link_in_slave_11_tready(link_in[11].slave.tReady),
        .link_in_master_12_tvalid(link_in[12].master.tValid),
        .link_in_master_12_tdata(link_in[12].master.tData),
        .link_in_master_12_tuser(link_in[12].master.tUser),
        .link_in_master_12_tlast(link_in[12].master.tLast),
        .link_in_slave_12_tready(link_in[12].slave.tReady),
        .link_in_master_13_tvalid(link_in[13].master.tValid),
        .link_in_master_13_tdata(link_in[13].master.tData),
        .link_in_master_13_tuser(link_in[13].master.tUser),
        .link_in_master_13_tlast(link_in[13].master.tLast),
        .link_in_slave_13_tready(link_in[13].slave.tReady),
        .link_in_master_14_tvalid(link_in[14].master.tValid),
        .link_in_master_14_tdata(link_in[14].master.tData),
        .link_in_master_14_tuser(link_in[14].master.tUser),
        .link_in_master_14_tlast(link_in[14].master.tLast),
        .link_in_slave_14_tready(link_in[14].slave.tReady),
        .link_in_master_15_tvalid(link_in[15].master.tValid),
        .link_in_master_15_tdata(link_in[15].master.tData),
        .link_in_master_15_tuser(link_in[15].master.tUser),
        .link_in_master_15_tlast(link_in[15].master.tLast),
        .link_in_slave_15_tready(link_in[15].slave.tReady),
        .link_in_master_16_tvalid(link_in[16].master.tValid),
        .link_in_master_16_tdata(link_in[16].master.tData),
        .link_in_master_16_tuser(link_in[16].master.tUser),
        .link_in_master_16_tlast(link_in[16].master.tLast),
        .link_in_slave_16_tready(link_in[16].slave.tReady),
        .link_in_master_17_tvalid(link_in[17].master.tValid),
        .link_in_master_17_tdata(link_in[17].master.tData),
        .link_in_master_17_tuser(link_in[17].master.tUser),
        .link_in_master_17_tlast(link_in[17].master.tLast),
        .link_in_slave_17_tready(link_in[17].slave.tReady),
        .link_in_master_18_tvalid(link_in[18].master.tValid),
        .link_in_master_18_tdata(link_in[18].master.tData),
        .link_in_master_18_tuser(link_in[18].master.tUser),
        .link_in_master_18_tlast(link_in[18].master.tLast),
        .link_in_slave_18_tready(link_in[18].slave.tReady),
        .link_in_master_19_tvalid(link_in[19].master.tValid),
        .link_in_master_19_tdata(link_in[19].master.tData),
        .link_in_master_19_tuser(link_in[19].master.tUser),
        .link_in_master_19_tlast(link_in[19].master.tLast),
        .link_in_slave_19_tready(link_in[19].slave.tReady),
        .link_in_master_20_tvalid(link_in[20].master.tValid),
        .link_in_master_20_tdata(link_in[20].master.tData),
        .link_in_master_20_tuser(link_in[20].master.tUser),
        .link_in_master_20_tlast(link_in[20].master.tLast),
        .link_in_slave_20_tready(link_in[20].slave.tReady),
        .link_in_master_21_tvalid(link_in[21].master.tValid),
        .link_in_master_21_tdata(link_in[21].master.tData),
        .link_in_master_21_tuser(link_in[21].master.tUser),
        .link_in_master_21_tlast(link_in[21].master.tLast),
        .link_in_slave_21_tready(link_in[21].slave.tReady),
        .link_in_master_22_tvalid(link_in[22].master.tValid),
        .link_in_master_22_tdata(link_in[22].master.tData),
        .link_in_master_22_tuser(link_in[22].master.tUser),
        .link_in_master_22_tlast(link_in[22].master.tLast),
        .link_in_slave_22_tready(link_in[22].slave.tReady),
        .link_in_master_23_tvalid(link_in[23].master.tValid),
        .link_in_master_23_tdata(link_in[23].master.tData),
        .link_in_master_23_tuser(link_in[23].master.tUser),
        .link_in_master_23_tlast(link_in[23].master.tLast),
        .link_in_slave_23_tready(link_in[23].slave.tReady),

        .link_out_master_0_tvalid(link_out[0].master.tValid),
        .link_out_master_0_tdata(link_out[0].master.tData),
        .link_out_master_0_tuser(link_out[0].master.tUser),
        .link_out_master_0_tlast(link_out[0].master.tLast),
        .link_out_slave_0_tready(link_out[0].slave.tReady),
        .link_out_master_1_tvalid(link_out[1].master.tValid),
        .link_out_master_1_tdata(link_out[1].master.tData),
        .link_out_master_1_tuser(link_out[1].master.tUser),
        .link_out_master_1_tlast(link_out[1].master.tLast),
        .link_out_slave_1_tready(link_out[1].slave.tReady),
        .link_out_master_2_tvalid(link_out[2].master.tValid),
        .link_out_master_2_tdata(link_out[2].master.tData),
        .link_out_master_2_tuser(link_out[2].master.tUser),
        .link_out_master_2_tlast(link_out[2].master.tLast),
        .link_out_slave_2_tready(link_out[2].slave.tReady),
        .link_out_master_3_tvalid(link_out[3].master.tValid),
        .link_out_master_3_tdata(link_out[3].master.tData),
        .link_out_master_3_tuser(link_out[3].master.tUser),
        .link_out_master_3_tlast(link_out[3].master.tLast),
        .link_out_slave_3_tready(link_out[3].slave.tReady),
        .link_out_master_4_tvalid(link_out[4].master.tValid),
        .link_out_master_4_tdata(link_out[4].master.tData),
        .link_out_master_4_tuser(link_out[4].master.tUser),
        .link_out_master_4_tlast(link_out[4].master.tLast),
        .link_out_slave_4_tready(link_out[4].slave.tReady),
        .link_out_master_5_tvalid(link_out[5].master.tValid),
        .link_out_master_5_tdata(link_out[5].master.tData),
        .link_out_master_5_tuser(link_out[5].master.tUser),
        .link_out_master_5_tlast(link_out[5].master.tLast),
        .link_out_slave_5_tready(link_out[5].slave.tReady),
        .link_out_master_6_tvalid(link_out[6].master.tValid),
        .link_out_master_6_tdata(link_out[6].master.tData),
        .link_out_master_6_tuser(link_out[6].master.tUser),
        .link_out_master_6_tlast(link_out[6].master.tLast),
        .link_out_slave_6_tready(link_out[6].slave.tReady),
        .link_out_master_7_tvalid(link_out[7].master.tValid),
        .link_out_master_7_tdata(link_out[7].master.tData),
        .link_out_master_7_tuser(link_out[7].master.tUser),
        .link_out_master_7_tlast(link_out[7].master.tLast),
        .link_out_slave_7_tready(link_out[7].slave.tReady),
        .link_out_master_8_tvalid(link_out[8].master.tValid),
        .link_out_master_8_tdata(link_out[8].master.tData),
        .link_out_master_8_tuser(link_out[8].master.tUser),
        .link_out_master_8_tlast(link_out[8].master.tLast),
        .link_out_slave_8_tready(link_out[8].slave.tReady),
        .link_out_master_9_tvalid(link_out[9].master.tValid),
        .link_out_master_9_tdata(link_out[9].master.tData),
        .link_out_master_9_tuser(link_out[9].master.tUser),
        .link_out_master_9_tlast(link_out[9].master.tLast),
        .link_out_slave_9_tready(link_out[9].slave.tReady),
        .link_out_master_10_tvalid(link_out[10].master.tValid),
        .link_out_master_10_tdata(link_out[10].master.tData),
        .link_out_master_10_tuser(link_out[10].master.tUser),
        .link_out_master_10_tlast(link_out[10].master.tLast),
        .link_out_slave_10_tready(link_out[10].slave.tReady),
        .link_out_master_11_tvalid(link_out[11].master.tValid),
        .link_out_master_11_tdata(link_out[11].master.tData),
        .link_out_master_11_tuser(link_out[11].master.tUser),
        .link_out_master_11_tlast(link_out[11].master.tLast),
        .link_out_slave_11_tready(link_out[11].slave.tReady),
        .link_out_master_12_tvalid(link_out[12].master.tValid),
        .link_out_master_12_tdata(link_out[12].master.tData),
        .link_out_master_12_tuser(link_out[12].master.tUser),
        .link_out_master_12_tlast(link_out[12].master.tLast),
        .link_out_slave_12_tready(link_out[12].slave.tReady),
        .link_out_master_13_tvalid(link_out[13].master.tValid),
        .link_out_master_13_tdata(link_out[13].master.tData),
        .link_out_master_13_tuser(link_out[13].master.tUser),
        .link_out_master_13_tlast(link_out[13].master.tLast),
        .link_out_slave_13_tready(link_out[13].slave.tReady),
        .link_out_master_14_tvalid(link_out[14].master.tValid),
        .link_out_master_14_tdata(link_out[14].master.tData),
        .link_out_master_14_tuser(link_out[14].master.tUser),
        .link_out_master_14_tlast(link_out[14].master.tLast),
        .link_out_slave_14_tready(link_out[14].slave.tReady),
        .link_out_master_15_tvalid(link_out[15].master.tValid),
        .link_out_master_15_tdata(link_out[15].master.tData),
        .link_out_master_15_tuser(link_out[15].master.tUser),
        .link_out_master_15_tlast(link_out[15].master.tLast),
        .link_out_slave_15_tready(link_out[15].slave.tReady),
        .link_out_master_16_tvalid(link_out[16].master.tValid),
        .link_out_master_16_tdata(link_out[16].master.tData),
        .link_out_master_16_tuser(link_out[16].master.tUser),
        .link_out_master_16_tlast(link_out[16].master.tLast),
        .link_out_slave_16_tready(link_out[16].slave.tReady),
        .link_out_master_17_tvalid(link_out[17].master.tValid),
        .link_out_master_17_tdata(link_out[17].master.tData),
        .link_out_master_17_tuser(link_out[17].master.tUser),
        .link_out_master_17_tlast(link_out[17].master.tLast),
        .link_out_slave_17_tready(link_out[17].slave.tReady),
        .link_out_master_18_tvalid(link_out[18].master.tValid),
        .link_out_master_18_tdata(link_out[18].master.tData),
        .link_out_master_18_tuser(link_out[18].master.tUser),
        .link_out_master_18_tlast(link_out[18].master.tLast),
        .link_out_slave_18_tready(link_out[18].slave.tReady),
        .link_out_master_19_tvalid(link_out[19].master.tValid),
        .link_out_master_19_tdata(link_out[19].master.tData),
        .link_out_master_19_tuser(link_out[19].master.tUser),
        .link_out_master_19_tlast(link_out[19].master.tLast),
        .link_out_slave_19_tready(link_out[19].slave.tReady),
        .link_out_master_20_tvalid(link_out[20].master.tValid),
        .link_out_master_20_tdata(link_out[20].master.tData),
        .link_out_master_20_tuser(link_out[20].master.tUser),
        .link_out_master_20_tlast(link_out[20].master.tLast),
        .link_out_slave_20_tready(link_out[20].slave.tReady),
        .link_out_master_21_tvalid(link_out[21].master.tValid),
        .link_out_master_21_tdata(link_out[21].master.tData),
        .link_out_master_21_tuser(link_out[21].master.tUser),
        .link_out_master_21_tlast(link_out[21].master.tLast),
        .link_out_slave_21_tready(link_out[21].slave.tReady),
        .link_out_master_22_tvalid(link_out[22].master.tValid),
        .link_out_master_22_tdata(link_out[22].master.tData),
        .link_out_master_22_tuser(link_out[22].master.tUser),
        .link_out_master_22_tlast(link_out[22].master.tLast),
        .link_out_slave_22_tready(link_out[22].slave.tReady),
        .link_out_master_23_tvalid(link_out[23].master.tValid),
        .link_out_master_23_tdata(link_out[23].master.tData),
        .link_out_master_23_tuser(link_out[23].master.tUser),
        .link_out_master_23_tlast(link_out[23].master.tLast),
        .link_out_slave_23_tready(link_out[23].slave.tReady)
    );


endmodule
