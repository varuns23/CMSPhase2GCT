library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

use work.StdRtlPkg.all;
use work.AxiStreamPkg.all;

entity algoStreamWrapper is
  generic (
    N_INPUT_STREAMS  : integer := 36;
    N_OUTPUT_STREAMS : integer := 36
    );
  port (
    -- Algo Control/Status Signals
    algoClk   : in  sl;
    algoRst   : in  sl;
    algoStart : in  sl;
    algoDone  : out sl := '0';
    algoIdle  : out sl := '0';
    algoReady : out sl := '0';

    -- AXI-Stream In/Out Ports
    axiStreamIn  : in  AxiStreamMasterArray(0 to N_INPUT_STREAMS-1);
    axiStreamOut : out AxiStreamMasterArray(0 to N_OUTPUT_STREAMS-1) := (others => AXI_STREAM_MASTER_INIT_C)
    );
end algoStreamWrapper;

architecture rtl of algoStreamWrapper is

  signal algoRstD1, algoRstD1n : sl;
  signal algoStartD1           : sl;

begin

  algoRstD1  <= algoRst when rising_edge(algoClk);
  algoRstD1n <= not algoRstD1;

  algoStartD1 <= algoStart when rising_edge(algoClk);

  U_algoStream : entity work.algoStream
    port map (
      ap_clk   => algoClk,
      ap_rst_n => algoRstD1n,
      ap_start => algoStartD1,
      ap_done  => algoDone,
      ap_idle  => algoIdle,
      ap_ready => algoReady,

      link_in_0_TUSER      => axiStreamIn(0).tUser(7 downto 0),
      link_in_0_TDATA      => axiStreamIn(0).tData(63 downto 0),
      link_in_0_TVALID     => axiStreamIn(0).tValid,
      link_in_0_TLAST(0)   => axiStreamIn(0).tLast,
      link_in_0_TREADY     => open,
      link_in_1_TUSER      => axiStreamIn(1).tUser(7 downto 0),
      link_in_1_TDATA      => axiStreamIn(1).tData(63 downto 0),
      link_in_1_TVALID     => axiStreamIn(1).tValid,
      link_in_1_TLAST(0)   => axiStreamIn(1).tLast,
      link_in_1_TREADY     => open,
      link_in_2_TUSER      => axiStreamIn(2).tUser(7 downto 0),
      link_in_2_TDATA      => axiStreamIn(2).tData(63 downto 0),
      link_in_2_TVALID     => axiStreamIn(2).tValid,
      link_in_2_TLAST(0)   => axiStreamIn(2).tLast,
      link_in_2_TREADY     => open,
      link_in_3_TUSER      => axiStreamIn(3).tUser(7 downto 0),
      link_in_3_TDATA      => axiStreamIn(3).tData(63 downto 0),
      link_in_3_TVALID     => axiStreamIn(3).tValid,
      link_in_3_TLAST(0)   => axiStreamIn(3).tLast,
      link_in_3_TREADY     => open,
      link_in_4_TUSER      => axiStreamIn(4).tUser(7 downto 0),
      link_in_4_TDATA      => axiStreamIn(4).tData(63 downto 0),
      link_in_4_TVALID     => axiStreamIn(4).tValid,
      link_in_4_TLAST(0)   => axiStreamIn(4).tLast,
      link_in_4_TREADY     => open,
      link_in_5_TUSER      => axiStreamIn(5).tUser(7 downto 0),
      link_in_5_TDATA      => axiStreamIn(5).tData(63 downto 0),
      link_in_5_TVALID     => axiStreamIn(5).tValid,
      link_in_5_TLAST(0)   => axiStreamIn(5).tLast,
      link_in_5_TREADY     => open,
      link_in_6_TUSER      => axiStreamIn(6).tUser(7 downto 0),
      link_in_6_TDATA      => axiStreamIn(6).tData(63 downto 0),
      link_in_6_TVALID     => axiStreamIn(6).tValid,
      link_in_6_TLAST(0)   => axiStreamIn(6).tLast,
      link_in_6_TREADY     => open,
      link_in_7_TUSER      => axiStreamIn(7).tUser(7 downto 0),
      link_in_7_TDATA      => axiStreamIn(7).tData(63 downto 0),
      link_in_7_TVALID     => axiStreamIn(7).tValid,
      link_in_7_TLAST(0)   => axiStreamIn(7).tLast,
      link_in_7_TREADY     => open,
      link_in_8_TUSER      => axiStreamIn(8).tUser(7 downto 0),
      link_in_8_TDATA      => axiStreamIn(8).tData(63 downto 0),
      link_in_8_TVALID     => axiStreamIn(8).tValid,
      link_in_8_TLAST(0)   => axiStreamIn(8).tLast,
      link_in_8_TREADY     => open,
      link_in_9_TUSER      => axiStreamIn(9).tUser(7 downto 0),
      link_in_9_TDATA      => axiStreamIn(9).tData(63 downto 0),
      link_in_9_TVALID     => axiStreamIn(9).tValid,
      link_in_9_TLAST(0)   => axiStreamIn(9).tLast,
      link_in_9_TREADY     => open,
      link_in_10_TUSER     => axiStreamIn(10).tUser(7 downto 0),
      link_in_10_TDATA     => axiStreamIn(10).tData(63 downto 0),
      link_in_10_TVALID    => axiStreamIn(10).tValid,
      link_in_10_TLAST(0)  => axiStreamIn(10).tLast,
      link_in_10_TREADY    => open,
      link_in_11_TUSER     => axiStreamIn(11).tUser(7 downto 0),
      link_in_11_TDATA     => axiStreamIn(11).tData(63 downto 0),
      link_in_11_TVALID    => axiStreamIn(11).tValid,
      link_in_11_TLAST(0)  => axiStreamIn(11).tLast,
      link_in_11_TREADY    => open,
      link_in_12_TUSER     => axiStreamIn(12).tUser(7 downto 0),
      link_in_12_TDATA     => axiStreamIn(12).tData(63 downto 0),
      link_in_12_TVALID    => axiStreamIn(12).tValid,
      link_in_12_TLAST(0)  => axiStreamIn(12).tLast,
      link_in_12_TREADY    => open,
      link_in_13_TUSER     => axiStreamIn(13).tUser(7 downto 0),
      link_in_13_TDATA     => axiStreamIn(13).tData(63 downto 0),
      link_in_13_TVALID    => axiStreamIn(13).tValid,
      link_in_13_TLAST(0)  => axiStreamIn(13).tLast,
      link_in_13_TREADY    => open,
      link_in_14_TUSER     => axiStreamIn(14).tUser(7 downto 0),
      link_in_14_TDATA     => axiStreamIn(14).tData(63 downto 0),
      link_in_14_TVALID    => axiStreamIn(14).tValid,
      link_in_14_TLAST(0)  => axiStreamIn(14).tLast,
      link_in_14_TREADY    => open,
      link_in_15_TUSER     => axiStreamIn(15).tUser(7 downto 0),
      link_in_15_TDATA     => axiStreamIn(15).tData(63 downto 0),
      link_in_15_TVALID    => axiStreamIn(15).tValid,
      link_in_15_TLAST(0)  => axiStreamIn(15).tLast,
      link_in_15_TREADY    => open,
      link_in_16_TUSER     => axiStreamIn(16).tUser(7 downto 0),
      link_in_16_TDATA     => axiStreamIn(16).tData(63 downto 0),
      link_in_16_TVALID    => axiStreamIn(16).tValid,
      link_in_16_TLAST(0)  => axiStreamIn(16).tLast,
      link_in_16_TREADY    => open,
      link_in_17_TUSER     => axiStreamIn(17).tUser(7 downto 0),
      link_in_17_TDATA     => axiStreamIn(17).tData(63 downto 0),
      link_in_17_TVALID    => axiStreamIn(17).tValid,
      link_in_17_TLAST(0)  => axiStreamIn(17).tLast,
      link_in_17_TREADY    => open,
      link_in_18_TUSER     => axiStreamIn(18).tUser(7 downto 0),
      link_in_18_TDATA     => axiStreamIn(18).tData(63 downto 0),
      link_in_18_TVALID    => axiStreamIn(18).tValid,
      link_in_18_TLAST(0)  => axiStreamIn(18).tLast,
      link_in_18_TREADY    => open,
      link_in_19_TUSER     => axiStreamIn(19).tUser(7 downto 0),
      link_in_19_TDATA     => axiStreamIn(19).tData(63 downto 0),
      link_in_19_TVALID    => axiStreamIn(19).tValid,
      link_in_19_TLAST(0)  => axiStreamIn(19).tLast,
      link_in_19_TREADY    => open,
      link_in_20_TUSER     => axiStreamIn(20).tUser(7 downto 0),
      link_in_20_TDATA     => axiStreamIn(20).tData(63 downto 0),
      link_in_20_TVALID    => axiStreamIn(20).tValid,
      link_in_20_TLAST(0)  => axiStreamIn(20).tLast,
      link_in_20_TREADY    => open, 
      link_in_21_TUSER     => axiStreamIn(21).tUser(7 downto 0),
      link_in_21_TDATA     => axiStreamIn(21).tData(63 downto 0),
      link_in_21_TVALID    => axiStreamIn(21).tValid,
      link_in_21_TLAST(0)  => axiStreamIn(21).tLast,
      link_in_21_TREADY    => open, 
      link_in_22_TUSER     => axiStreamIn(22).tUser(7 downto 0),
      link_in_22_TDATA     => axiStreamIn(22).tData(63 downto 0),
      link_in_22_TVALID    => axiStreamIn(22).tValid,
      link_in_22_TLAST(0)  => axiStreamIn(22).tLast,
      link_in_22_TREADY    => open, 
      link_in_23_TUSER     => axiStreamIn(23).tUser(7 downto 0),
      link_in_23_TDATA     => axiStreamIn(23).tData(63 downto 0),
      link_in_23_TVALID    => axiStreamIn(23).tValid,
      link_in_23_TLAST(0)  => axiStreamIn(23).tLast,
      link_in_23_TREADY    => open, 
      link_in_24_TUSER     => axiStreamIn(24).tUser(7 downto 0),
      link_in_24_TDATA     => axiStreamIn(24).tData(63 downto 0),
      link_in_24_TVALID    => axiStreamIn(24).tValid,
      link_in_24_TLAST(0)  => axiStreamIn(24).tLast,
      link_in_24_TREADY    => open, 
      link_in_25_TUSER     => axiStreamIn(25).tUser(7 downto 0),
      link_in_25_TDATA     => axiStreamIn(25).tData(63 downto 0),
      link_in_25_TVALID    => axiStreamIn(25).tValid,
      link_in_25_TLAST(0)  => axiStreamIn(25).tLast,
      link_in_25_TREADY    => open, 
      link_in_26_TUSER     => axiStreamIn(26).tUser(7 downto 0),
      link_in_26_TDATA     => axiStreamIn(26).tData(63 downto 0),
      link_in_26_TVALID    => axiStreamIn(26).tValid,
      link_in_26_TLAST(0)  => axiStreamIn(26).tLast,
      link_in_26_TREADY    => open, 
      link_in_27_TUSER     => axiStreamIn(27).tUser(7 downto 0),
      link_in_27_TDATA     => axiStreamIn(27).tData(63 downto 0),
      link_in_27_TVALID    => axiStreamIn(27).tValid,
      link_in_27_TLAST(0)  => axiStreamIn(27).tLast,
      link_in_27_TREADY    => open, 
      link_in_28_TUSER     => axiStreamIn(28).tUser(7 downto 0),
      link_in_28_TDATA     => axiStreamIn(28).tData(63 downto 0),
      link_in_28_TVALID    => axiStreamIn(28).tValid,
      link_in_28_TLAST(0)  => axiStreamIn(28).tLast,
      link_in_28_TREADY    => open, 
      link_in_29_TUSER     => axiStreamIn(29).tUser(7 downto 0),
      link_in_29_TDATA     => axiStreamIn(29).tData(63 downto 0),
      link_in_29_TVALID    => axiStreamIn(29).tValid,
      link_in_29_TLAST(0)  => axiStreamIn(29).tLast,
      link_in_29_TREADY    => open, 
      link_in_30_TUSER     => axiStreamIn(30).tUser(7 downto 0),
      link_in_30_TDATA     => axiStreamIn(30).tData(63 downto 0),
      link_in_30_TVALID    => axiStreamIn(30).tValid,
      link_in_30_TLAST(0)  => axiStreamIn(30).tLast,
      link_in_30_TREADY    => open, 
      link_in_31_TUSER     => axiStreamIn(31).tUser(7 downto 0),
      link_in_31_TDATA     => axiStreamIn(31).tData(63 downto 0),
      link_in_31_TVALID    => axiStreamIn(31).tValid,
      link_in_31_TLAST(0)  => axiStreamIn(31).tLast,
      link_in_31_TREADY    => open, 
      link_in_32_TUSER     => axiStreamIn(32).tUser(7 downto 0),
      link_in_32_TDATA     => axiStreamIn(32).tData(63 downto 0),
      link_in_32_TVALID    => axiStreamIn(32).tValid,
      link_in_32_TLAST(0)  => axiStreamIn(32).tLast,
      link_in_32_TREADY    => open, 
      link_in_33_TUSER     => axiStreamIn(33).tUser(7 downto 0),
      link_in_33_TDATA     => axiStreamIn(33).tData(63 downto 0),
      link_in_33_TVALID    => axiStreamIn(33).tValid,
      link_in_33_TLAST(0)  => axiStreamIn(33).tLast,
      link_in_33_TREADY    => open, 
      link_in_34_TUSER     => axiStreamIn(34).tUser(7 downto 0),
      link_in_34_TDATA     => axiStreamIn(34).tData(63 downto 0),
      link_in_34_TVALID    => axiStreamIn(34).tValid,
      link_in_34_TLAST(0)  => axiStreamIn(34).tLast,
      link_in_34_TREADY    => open, 
      link_in_35_TUSER     => axiStreamIn(35).tUser(7 downto 0),
      link_in_35_TDATA     => axiStreamIn(35).tData(63 downto 0),
      link_in_35_TVALID    => axiStreamIn(35).tValid,
      link_in_35_TLAST(0)  => axiStreamIn(35).tLast,
      link_in_35_TREADY    => open, 
      link_out_0_TUSER     => axiStreamOut(0).tUser(7 downto 0),
      link_out_0_TDATA     => axiStreamOut(0).tData(63 downto 0),
      link_out_0_TVALID    => axiStreamOut(0).tValid,
      link_out_0_TLAST(0)  => axiStreamOut(0).tLast,
      link_out_0_TREADY    => '1', 
      link_out_1_TUSER     => axiStreamOut(1).tUser(7 downto 0),
      link_out_1_TDATA     => axiStreamOut(1).tData(63 downto 0),
      link_out_1_TVALID    => axiStreamOut(1).tValid,
      link_out_1_TLAST(0)  => axiStreamOut(1).tLast,
      link_out_1_TREADY    => '1', 
      link_out_2_TUSER     => axiStreamOut(2).tUser(7 downto 0),
      link_out_2_TDATA     => axiStreamOut(2).tData(63 downto 0),
      link_out_2_TVALID    => axiStreamOut(2).tValid,
      link_out_2_TLAST(0)  => axiStreamOut(2).tLast,
      link_out_2_TREADY    => '1', 
      link_out_3_TUSER     => axiStreamOut(3).tUser(7 downto 0),
      link_out_3_TDATA     => axiStreamOut(3).tData(63 downto 0),
      link_out_3_TVALID    => axiStreamOut(3).tValid,
      link_out_3_TLAST(0)  => axiStreamOut(3).tLast,
      link_out_3_TREADY    => '1', 
      link_out_4_TUSER     => axiStreamOut(4).tUser(7 downto 0),
      link_out_4_TDATA     => axiStreamOut(4).tData(63 downto 0),
      link_out_4_TVALID    => axiStreamOut(4).tValid,
      link_out_4_TLAST(0)  => axiStreamOut(4).tLast,
      link_out_4_TREADY    => '1', 
      link_out_5_TUSER     => axiStreamOut(5).tUser(7 downto 0),
      link_out_5_TDATA     => axiStreamOut(5).tData(63 downto 0),
      link_out_5_TVALID    => axiStreamOut(5).tValid,
      link_out_5_TLAST(0)  => axiStreamOut(5).tLast,
      link_out_5_TREADY    => '1', 
      link_out_6_TUSER     => axiStreamOut(6).tUser(7 downto 0),
      link_out_6_TDATA     => axiStreamOut(6).tData(63 downto 0),
      link_out_6_TVALID    => axiStreamOut(6).tValid,
      link_out_6_TLAST(0)  => axiStreamOut(6).tLast,
      link_out_6_TREADY    => '1', 
      link_out_7_TUSER     => axiStreamOut(7).tUser(7 downto 0),
      link_out_7_TDATA     => axiStreamOut(7).tData(63 downto 0),
      link_out_7_TVALID    => axiStreamOut(7).tValid,
      link_out_7_TLAST(0)  => axiStreamOut(7).tLast,
      link_out_7_TREADY    => '1', 
      link_out_8_TUSER     => axiStreamOut(8).tUser(7 downto 0),
      link_out_8_TDATA     => axiStreamOut(8).tData(63 downto 0),
      link_out_8_TVALID    => axiStreamOut(8).tValid,
      link_out_8_TLAST(0)  => axiStreamOut(8).tLast,
      link_out_8_TREADY    => '1', 
      link_out_9_TUSER     => axiStreamOut(9).tUser(7 downto 0),
      link_out_9_TDATA     => axiStreamOut(9).tData(63 downto 0),
      link_out_9_TVALID    => axiStreamOut(9).tValid,
      link_out_9_TLAST(0)  => axiStreamOut(9).tLast,
      link_out_9_TREADY    => '1', 
      link_out_10_TUSER    => axiStreamOut(10).tUser(7 downto 0),
      link_out_10_TDATA    => axiStreamOut(10).tData(63 downto 0),
      link_out_10_TVALID   => axiStreamOut(10).tValid,
      link_out_10_TLAST(0) => axiStreamOut(10).tLast,
      link_out_10_TREADY   => '1', 
      link_out_11_TUSER    => axiStreamOut(11).tUser(7 downto 0),
      link_out_11_TDATA    => axiStreamOut(11).tData(63 downto 0),
      link_out_11_TVALID   => axiStreamOut(11).tValid,
      link_out_11_TLAST(0) => axiStreamOut(11).tLast,
      link_out_11_TREADY   => '1', 
      link_out_12_TUSER    => axiStreamOut(12).tUser(7 downto 0),
      link_out_12_TDATA    => axiStreamOut(12).tData(63 downto 0),
      link_out_12_TVALID   => axiStreamOut(12).tValid,
      link_out_12_TLAST(0) => axiStreamOut(12).tLast,
      link_out_12_TREADY   => '1', 
      link_out_13_TUSER    => axiStreamOut(13).tUser(7 downto 0),
      link_out_13_TDATA    => axiStreamOut(13).tData(63 downto 0),
      link_out_13_TVALID   => axiStreamOut(13).tValid,
      link_out_13_TLAST(0) => axiStreamOut(13).tLast,
      link_out_13_TREADY   => '1', 
      link_out_14_TUSER    => axiStreamOut(14).tUser(7 downto 0),
      link_out_14_TDATA    => axiStreamOut(14).tData(63 downto 0),
      link_out_14_TVALID   => axiStreamOut(14).tValid,
      link_out_14_TLAST(0) => axiStreamOut(14).tLast,
      link_out_14_TREADY   => '1', 
      link_out_15_TUSER    => axiStreamOut(15).tUser(7 downto 0),
      link_out_15_TDATA    => axiStreamOut(15).tData(63 downto 0),
      link_out_15_TVALID   => axiStreamOut(15).tValid,
      link_out_15_TLAST(0) => axiStreamOut(15).tLast,
      link_out_15_TREADY   => '1', 
      link_out_16_TUSER    => axiStreamOut(16).tUser(7 downto 0),
      link_out_16_TDATA    => axiStreamOut(16).tData(63 downto 0),
      link_out_16_TVALID   => axiStreamOut(16).tValid,
      link_out_16_TLAST(0) => axiStreamOut(16).tLast,
      link_out_16_TREADY   => '1', 
      link_out_17_TUSER    => axiStreamOut(17).tUser(7 downto 0),
      link_out_17_TDATA    => axiStreamOut(17).tData(63 downto 0),
      link_out_17_TVALID   => axiStreamOut(17).tValid,
      link_out_17_TLAST(0) => axiStreamOut(17).tLast,
      link_out_17_TREADY   => '1', 
      link_out_18_TUSER    => axiStreamOut(18).tUser(7 downto 0),
      link_out_18_TDATA    => axiStreamOut(18).tData(63 downto 0),
      link_out_18_TVALID   => axiStreamOut(18).tValid,
      link_out_18_TLAST(0) => axiStreamOut(18).tLast,
      link_out_18_TREADY   => '1', 
      link_out_19_TUSER    => axiStreamOut(19).tUser(7 downto 0),
      link_out_19_TDATA    => axiStreamOut(19).tData(63 downto 0),
      link_out_19_TVALID   => axiStreamOut(19).tValid,
      link_out_19_TLAST(0) => axiStreamOut(19).tLast,
      link_out_19_TREADY   => '1', 
      link_out_20_TUSER    => axiStreamOut(20).tUser(7 downto 0),
      link_out_20_TDATA    => axiStreamOut(20).tData(63 downto 0),
      link_out_20_TVALID   => axiStreamOut(20).tValid,
      link_out_20_TLAST(0) => axiStreamOut(20).tLast,
      link_out_20_TREADY   => '1', 
      link_out_21_TUSER    => axiStreamOut(21).tUser(7 downto 0),
      link_out_21_TDATA    => axiStreamOut(21).tData(63 downto 0),
      link_out_21_TVALID   => axiStreamOut(21).tValid,
      link_out_21_TLAST(0) => axiStreamOut(21).tLast,
      link_out_21_TREADY   => '1', 
      link_out_22_TUSER    => axiStreamOut(22).tUser(7 downto 0),
      link_out_22_TDATA    => axiStreamOut(22).tData(63 downto 0),
      link_out_22_TVALID   => axiStreamOut(22).tValid,
      link_out_22_TLAST(0) => axiStreamOut(22).tLast,
      link_out_22_TREADY   => '1', 
      link_out_23_TUSER    => axiStreamOut(23).tUser(7 downto 0),
      link_out_23_TDATA    => axiStreamOut(23).tData(63 downto 0),
      link_out_23_TVALID   => axiStreamOut(23).tValid,
      link_out_23_TLAST(0) => axiStreamOut(23).tLast,
      link_out_23_TREADY   => '1', 
      link_out_24_TUSER    => axiStreamOut(24).tUser(7 downto 0),
      link_out_24_TDATA    => axiStreamOut(24).tData(63 downto 0),
      link_out_24_TVALID   => axiStreamOut(24).tValid,
      link_out_24_TLAST(0) => axiStreamOut(24).tLast,
      link_out_24_TREADY   => '1', 
      link_out_25_TUSER    => axiStreamOut(25).tUser(7 downto 0),
      link_out_25_TDATA    => axiStreamOut(25).tData(63 downto 0),
      link_out_25_TVALID   => axiStreamOut(25).tValid,
      link_out_25_TLAST(0) => axiStreamOut(25).tLast,
      link_out_25_TREADY   => '1', 
      link_out_26_TUSER    => axiStreamOut(26).tUser(7 downto 0),
      link_out_26_TDATA    => axiStreamOut(26).tData(63 downto 0),
      link_out_26_TVALID   => axiStreamOut(26).tValid,
      link_out_26_TLAST(0) => axiStreamOut(26).tLast,
      link_out_26_TREADY   => '1', 
      link_out_27_TUSER    => axiStreamOut(27).tUser(7 downto 0),
      link_out_27_TDATA    => axiStreamOut(27).tData(63 downto 0),
      link_out_27_TVALID   => axiStreamOut(27).tValid,
      link_out_27_TLAST(0) => axiStreamOut(27).tLast,
      link_out_27_TREADY   => '1', 
      link_out_28_TUSER    => axiStreamOut(28).tUser(7 downto 0),
      link_out_28_TDATA    => axiStreamOut(28).tData(63 downto 0),
      link_out_28_TVALID   => axiStreamOut(28).tValid,
      link_out_28_TLAST(0) => axiStreamOut(28).tLast,
      link_out_28_TREADY   => '1', 
      link_out_29_TUSER    => axiStreamOut(29).tUser(7 downto 0),
      link_out_29_TDATA    => axiStreamOut(29).tData(63 downto 0),
      link_out_29_TVALID   => axiStreamOut(29).tValid,
      link_out_29_TLAST(0) => axiStreamOut(29).tLast,
      link_out_29_TREADY   => '1', 
      link_out_30_TUSER    => axiStreamOut(30).tUser(7 downto 0),
      link_out_30_TDATA    => axiStreamOut(30).tData(63 downto 0),
      link_out_30_TVALID   => axiStreamOut(30).tValid,
      link_out_30_TLAST(0) => axiStreamOut(30).tLast,
      link_out_30_TREADY   => '1', 
      link_out_31_TUSER    => axiStreamOut(31).tUser(7 downto 0),
      link_out_31_TDATA    => axiStreamOut(31).tData(63 downto 0),
      link_out_31_TVALID   => axiStreamOut(31).tValid,
      link_out_31_TLAST(0) => axiStreamOut(31).tLast,
      link_out_31_TREADY   => '1', 
      link_out_32_TUSER    => axiStreamOut(32).tUser(7 downto 0),
      link_out_32_TDATA    => axiStreamOut(32).tData(63 downto 0),
      link_out_32_TVALID   => axiStreamOut(32).tValid,
      link_out_32_TLAST(0) => axiStreamOut(32).tLast,
      link_out_32_TREADY   => '1', 
      link_out_33_TUSER    => axiStreamOut(33).tUser(7 downto 0),
      link_out_33_TDATA    => axiStreamOut(33).tData(63 downto 0),
      link_out_33_TVALID   => axiStreamOut(33).tValid,
      link_out_33_TLAST(0) => axiStreamOut(33).tLast,
      link_out_33_TREADY   => '1', 
      link_out_34_TUSER    => axiStreamOut(34).tUser(7 downto 0),
      link_out_34_TDATA    => axiStreamOut(34).tData(63 downto 0),
      link_out_34_TVALID   => axiStreamOut(34).tValid,
      link_out_34_TLAST(0) => axiStreamOut(34).tLast,
      link_out_34_TREADY   => '1', 
      link_out_35_TUSER    => axiStreamOut(35).tUser(7 downto 0),
      link_out_35_TDATA    => axiStreamOut(35).tData(63 downto 0),
      link_out_35_TVALID   => axiStreamOut(35).tValid,
      link_out_35_TLAST(0) => axiStreamOut(35).tLast,
      link_out_35_TREADY   => '1' 
      );


end rtl;
